# ====================================================================
#
#      i2c_mips_vcoreiii.cdl
#
#      eCos mips VCOREIIII2C configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2005, 2006 eCosCentric Limited
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Lars Povlsen
# Contributors:   
# Date:           2010-08-04
#
#####DESCRIPTIONEND####
# ====================================================================


cdl_package CYGPKG_IO_I2C_MIPS_VCOREIII {
    display         "I2C driver for Vitesse Semiconductior VCOREIII family"

    parent          CYGPKG_IO_I2C
    active_if       CYGPKG_IO_I2C
    active_if       CYGPKG_IO_I2C
	
    description   "
           This package provides a generic I2C device driver for the on-chip
           I2C modules in Vitesse VCOREIII processors."

    include_dir     cyg/io
    compile 	    i2c_vcoreiii.c

    cdl_component CYGPKG_DEVS_I2C_VCOREIII_OPTIONS {
        display 	"I2C driver build options"
        flavor  	none
	active_if	{ CYGINT_DEVS_I2C_VCOREIII_BUS_DEVICES > 0 }
        description   "
	    Package specific build options including control over
	    compiler flags used only in building the VCOREIII I2C
            bus driver."

        cdl_option CYGPKG_DEVS_I2C_VCOREIII_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the VCOREIII I2C bus driver. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_I2C_VCOREIII_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the VCOREIII I2C bus driver. These flags are
                removed from the set of global flags if present."
        }
    }
}
