##=============================================================================
##
##      spi_vcoreiii.cdl
##
##      VCore-III SPI driver configuration options.
##
##=============================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##=============================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):       Lars Povlsen
## Contributors(s): Chris Holgate (based on CortexM STM32 code)
## Date:            2009-09-14
## Purpose:         Configure VCore-III SPI driver.
##
######DESCRIPTIONEND####
##
##=============================================================================

cdl_package CYGPKG_DEVS_SPI_MIPS_VCOREIII {
    display       "Vitesse VCore-III SPI driver"
    description   "
        This package provides SPI driver support for the Vitesse VCore-III processor
        family.
    "
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    requires      CYGPKG_HAL_MIPS_VCOREIII || CYGPKG_HAL_MIPS_VCOREIII_SERVAL
    hardware
    include_dir   cyg/io
    compile       spi_vcoreiii.c

    cdl_option CYGPKG_DEVS_SPI_MIPS_VCOREIII_TESTS {
            display "VCore-III SPI tests"
            flavor  data
            no_define
            calculated { "tests/spi1test" }
            description   "
                This option specifies the set of tests for the VCore-III SPI device driver."
    }

}
# EOF spi_vcoreiii.cdl
