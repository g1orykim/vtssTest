# ====================================================================
#
#      httpd.cdl
#
#      HTTP server configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2005 eCosCentric Ltd.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Anthony Tonizzo (atonizzo@gmail.com)
# Contributors:   
# Date:           2006-06-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_ATHTTPD {
    display       "Another Tiny HTTP server"
    description   "This package provides a small footprint web server for eCos
                   with configurable features."
    include_dir   cyg/athttpd
    include_files auth.h digcalc.h forms.h global.h handler.h http.h md5.h socket.h cgi.h jim.h
    compile       forms.c handler.c http.c socket.c cgi.c
    requires      CYGPKG_NET
    requires      !CYGPKG_HTTPD
# ====================================================================
   
    cdl_component CYGPKG_NET_ATHTTPD_THREADOPT {
        display "Thread settings"
        flavor  none
        no_define
        description   "Options to change certain thread values."

      cdl_option CYGNUM_NET_ATHTTPD_THREADOPT_PRIORITY {
          display "Thread priority"
          flavor data
          default_value { CYGNUM_KERNEL_SCHED_PRIORITIES/2 }
          legal_values 0 to CYGNUM_KERNEL_SCHED_PRIORITIES
          description "The HTTP server threads can be run at any priority.
                       The exact priority depends on the importance of the
                       server relative to the rest of the system. The default
                       is to put it in the middle of the priority range to provide
                       reasonable response without impacting genuine high
                       priority threads."
      }

      cdl_option CYGNUM_NET_ATHTTPD_THREADOPT_STACKSIZE {
          display "Thread stack size"
          flavor data
          default_value 4096
          description "This is the amount of extra stack to be allocated for 
                       the HTTPD thread. This value is added to
                       CYGNUM_HAL_STACK_SIZE_MINIMUM to determine the final
                       size of the stack for the server."
      }
    }  

    cdl_component CYGOPT_NET_ATHTTPD_SERVEROPT {
        display "Server settings"
        flavor  none
        no_define
        description   "Options to change certain server options."

      cdl_option CYGNUM_NET_ATHTTPD_SERVEROPT_PORT {
          display "Server Port"
          flavor data
          default_value 80
          description "This is the port on which the server will be listening
                      for requests. Unless overridden in the request by the 
                      client, the well known port for HTTP is 80."
      }

      cdl_option CYGDAT_NET_ATHTTPD_SERVEROPT_SERVERID {
          display "Server ID string"
          flavor data
          default_value {"\"eCos Embedded Web Server\""}
          description "This is the string sent out in the 'Server:' header line."
      }
      
      cdl_option CYGNUM_ATHTTPD_SERVER_BUFFER_SIZE {
          display "IO buffer size"
          flavor data
          default_value 10240
          description "This option defines the size of the buffers used to 
                       receive and transmit transmit data to and from the TCP/IP
                       stack.
                       The limit is in MSIE and Safari about 2KB, in Opera about
                       4KB and in Firefox about 8KB. We may thus assume that 8KB
                       is the maximum possible length and that 2KB is a more
                       affordable length to rely on at the server side and that
                       255 bytes is the safest length to assume that the entire
                       URL will come in."
      }

      cdl_option CYGNUM_ATHTTPD_SERVER_MAX_POST {
          display "Maximum data received upon POST"
          flavor data
          default_value 2048
          description "This option defines the size of maximum amount of data 
                       the web server will accept from POST'ed forms."
      }

      cdl_option CYGDAT_NET_ATHTTPD_SERVEROPT_ROOTDIR {
          display "HTTPD root directory"
          flavor data
          default_value {"\"/\""}
          description "This is the absolute path in the eCos file system to the 
                       HTML documents, including cgi-bin files and error
                       files and it is generally where the web server will
                       look for the index file. Include a trailing slash."
      }
      
      cdl_option CYGDAT_NET_ATHTTPD_SERVEROPT_CGIDIR {
          display "cgi-bin directory"
          active_if    { 0 != CYGOPT_NET_ATHTTPD_USE_CGIBIN_OBJLOADER || 0 != CYGOPT_NET_ATHTTPD_USE_CGIBIN_TCL }
          flavor data
          default_value {"\"cgi-bin/\""}
          description "This is the path, relative to CYGDAT_NET_ATHTTPD_SERVEROPT_ROOTDIR,
                       where the cgi-bin files are stored. Based on the extension
                       of the cgi-bin file requested, the appropriate interpreter
                       will be used. Include a trailing slash."
      }
      
      cdl_option CYGDAT_NET_ATHTTPD_SERVEROPT_ERRORDIR {
          display "Error files directory"
          flavor data
          default_value {"\"errors/\""}
          description "This is the path, relative to the CYGDAT_NET_ATHTTPD_SERVEROPT_ROOTDIR,
                       that contains the user-defined files that are sent out
                       by the server in case of error. The files are named
                       error_XXX.html where XXX is the 3 digit HTML code. 
                       For example, for a 404 error the server file will be
                       named error_404.html. Upon a 404 error, the server will
                       check the existence of such a file in this directory and
                       if found, it will send it out. Missing that file, a
                       standard simple message will be sent instead. Include 
                       a trailing slash."
      }

      cdl_option CYGDAT_NET_ATHTTPD_DEFAULT_MIME_TYPE {
          display "Default MIME type"
          flavor data
          default_value {"\"text/plain\""}
          description "When accessing internal resources or a file system,
                       the MIME type is determined by first finding the extension
                       of the file itself and then by looking up the extension
                       in the MIME table. In case no extension is found the user 
                       can define the default MIME type to use. Notice that
                       this is the full MIME type and not the extension.
                       A list of standard MIME types sorted by extension can
                       be found in the current/doc directory"
      }
      
      cdl_option CYGDAT_NET_ATHTTPD_ALTERNATE_HOME {
          display "User defined Home Page"
          flavor booldata
          default_value {"\"/index.html\""}
          description "This file name defines the name of a custom index file 
                       and is used in case none of the default index files are 
                       found in a directory. Notice that this file name is
                       only appended to GET requests for \"/\""
      }
    }  

    cdl_option CYGOPT_NET_ATHTTPD_USE_FS {
        display       "Support for file system access"
        flavor        bool
        default_value 1
        active_if     CYGPKG_IO_FILEIO
        description   "
            This option enables the use of a file system to access the pages
             to be served. It is the responsibility of the user to properly
             mount the file system(s) required by the web server. If this
             option is not selected each URL requested must be serviced using
             either c language callbacks or internal resources." 
    }

    cdl_option CYGOPT_NET_ATHTTPD_USE_AUTH {
        display       "Support for basic authentication"
        flavor        bool
        default_value 0
        description   "
            This option enables the use basic authentication in web pages.
            Digest authentication code is also included, but has not been
            extensively tested." 
       compile md5c.c
       compile auth.c
    }

    cdl_option CYGOPT_NET_ATHTTPD_BASIC_AUTH_MAX_USERNAME_LEN {
        display       "When using basic authentication, maximum length of user name"
        flavor        data
        default_value 32
        description   "
            This option defines the maximum length of the user name excluding
            terminating NULL, and is used only when CYGOPT_NET_ATHTTPD_USE_AUTH
            is enabled and the method is 'Basic'."
    }

    cdl_option CYGOPT_NET_ATHTTPD_BASIC_AUTH_MAX_PASSWORD_LEN {
        display       "When using basic authentication, maximum length of password"
        flavor        data
        default_value 32
        description   "
            This option defines the maximum length of the password excluding
            terminating NULL, and is used only when CYGOPT_NET_ATHTTPD_USE_AUTH
            is enabled and the method is 'Basic'."
    }

    cdl_option CYGOPT_NET_ATHTTPD_INIT_ALL_NETWORK_INTERFACES {
        display       "Call init_all_network_interfaces() when starting daemon?"
        flavor        bool
        default_value 1
        description   "
            Some applications may want to control the call to
            init_all_network_interfaces() themselves, for instance if
            using DHCP, and the application code wishes to control whether
            to start DHCP or not. Default is to call init_all_network_interfaces()."
    }

    cdl_option CYGOPT_NET_ATHTTPD_CLOSE_CHUNKED_CONNECTIONS {
        display       "Close connections used for chunked transfer"
        flavor        bool
        default_value 1
        description   "
            This option causes connections used for chunked transfer to be
             closed after use. Persisting the connection will use less
             network resources and will improve latency, but may do so at
             the risk of compatibility with older browsers."
    }

    cdl_option CYGOPT_NET_ATHTTPD_DOCUMENT_EXPIRATION_TIME {
        display          "Maximum lifetime of a document in seconds"
        flavor           data
        default_value    0
        description      "
            This options causes documents to 'expire' after a set number
            of seconds. If certain pages are updated frequently, it might be a
            good idea to assign them an expitation time in seconds. If the
            client needs to reload a page that has expired, it will request
            it again, otherwise it will use the copy in the cache. A value
            of 0 means that this option is disabled. Any other value
            represents the number of seconds (after the last modification to
            the document) after which the page becomes stale. This option
            applies to all the pages (including those that reside in ROM
            and thus, by definition, won't change) and thus is it preferable
            to use the CYG_HTTPD_MODE_NO_CACHE mode for pages that need to be
            refreshed frequently."
    }

    cdl_option CYGOPT_NET_ATHTTPD_HTTPS {
        display       "Support for HTTPS authentication."
        flavor        bool
        default_value 1
        description   "This option defines the HTTPS supported or not.
                       To enable the function, another eCos package 
                       CYGPKG_OPENSSL is required"
    }

    cdl_option CYGNUM_NET_ATHTTPD_HTTPS_SERVEROPT_PORT {
        display "HTTPS Server Port"
        flavor data
        default_value 443
        description "This is the port on which the HTTPS server will be listening
                    for requests. Unless overridden in the request by the 
                    client, the well known port for HTTP is 443."
    }

    cdl_option CYGOPT_NET_ATHTTPD_USE_DIRLIST {
        display       "Support for directory listing"
        flavor        bool
        default_value 0
        active_if     CYGPKG_IO_FILEIO
        active_if     CYGOPT_NET_ATHTTPD_USE_FS
        description   "
            When a client issues a request that ends in '/' the server will
            try to locate anyone of a number of index files. Failing to find
            one, it will list the directory contents."
    }

    cdl_component CYGOPT_NET_ATHTTPD_CGIBIN {
        display "Supported CGI Types"
        flavor  none
        no_define
        description   "Options to select which CGI types are supported."

      cdl_option CYGOPT_NET_ATHTTPD_USE_CGIBIN_OBJLOADER {
          display       "Support cgi via the OBJLOADER package"
          flavor        bool
          default_value 0
          active_if     CYGPKG_OBJLOADER
          description   "This option enables the use of the object loader 
                         package as a means of providing on-demand loading and 
                         execution of code, thus providing a simple cgi
                         capability that does not involve scripting." 
      }

      cdl_option CYGOPT_NET_ATHTTPD_USE_CGIBIN_TCL {
          display       "Support cgi via the a simple tcl interpreter (jim)"
          flavor        bool
          default_value 0
          description   "This option enables the use of a small tcl
                         interpreter as a means of providing a simple cgi
                         capability. Checking this option increases 
                         considerably the size of the executable." 
          compile       jim.c
          define        JIM_ANSIC
          define        JIM_EMBEDDED
      }
    }  

    cdl_option CYGOPT_NET_ATHTTPD_USE_IRES_ETAG {
        display       "Use ETag for client caching of internal ressources."
        flavor        bool
        default_value 0
        description   "
            This option causes internal resources to be made cacheable
            though the use of a 'extern char http_ires_etag[]' - which
            must be provide and initialized externally from
            ATHTTPD. Response headers for internal resources will
            include the ETag, and requests for internal resources
            will check whether a cached version is up to date (sending
            a '304 Not modified' response back)."

    }

    cdl_option CYGOPT_NET_ATHTTPD_USE_COOKIES {
        display       "Use HTTP cookies."
        flavor        bool
        default_value 0
        description   "
            This option causes internal resources to use HTTP cookie."
    }

    cdl_option CYGOPT_NET_ATHTTPD_USE_COOKIE_AUTH {
        display       "Use cookie to implement authentication."
        flavor        bool
        default_value 0
        description   "
            This option causes internal resources to use cookie instead
            of using HTTP basic authentication. The chief advantage of
            cookies is flexibility: we can handle the whole process ourself."
    }

    cdl_option CYGOPT_NET_ATHTTPD_USE_IRES_HEADER {
        display       "Use this HTTP header for all internal ressources"
        flavor        booldata
        default_value 0
        description   "
            This option defines a HTTP header sent for all internal
            resources. The header must end with a \\r\\n.
            Commonly, this can be used to control client-side caching."
    }

    cdl_option CYGOPT_NET_ATHTTPD_DEBUG_LEVEL {
        display          "Verbosity of debug output"
        flavor           data
        legal_values     0 1 2
        default_value    0
        description      "This option allows controls over the verbosity of
                         the debug output. 1 mostly reports opening and
                         closing of socket descriptors, 2 is very
                         verbose, including the name of all files sent
                         out, including internal resources."
    }
    cdl_component CYGPKG_ATHTTPD_OPTIONS {
        display "AT HTTP server build options"
        flavor  none
        no_define

        cdl_option CYGPKG_ATHTTPD_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the HTTP server package.
                These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_ATHTTPD_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the HTTP server package. These flags are removed from
                the set of global flags if present."
        }
    }
}

# ====================================================================
# EOF httpd.cdl
